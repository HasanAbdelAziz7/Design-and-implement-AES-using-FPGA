package AES_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"


`include"AES_sequencer.sv"
`include"AES_driver.sv"
`include"AES_monitor.sv"
`include"AES_agent.sv"
`include"AES_scoreboard.sv"
`include"AES_env.sv"
`include"AES_test.sv"

endpackage
